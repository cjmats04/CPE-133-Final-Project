`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: Cal Poly
// Engineer: Calvin Matsushita
// 
// Create Date: 
// Design Name: 
// Module Name: 
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module TK_TB();

	logic clk;
	logic TB_EN;
	logic TB_RST;
	logic [3:0] TB_A;
	logic [3:0] TB_B;
	logic TB_P1L;
	logic TB_P2L;
	logic TB_CLR;

	TK UUT(.clk(clk), .TK_EN(TB_EN), .TK_RST(TB_RST), .TK_A(TB_A), .TK_B(TB_B), .TK_P1L(TB_P1L), .TK_P2L(TB_P2L), .TK_CLR(TB_CLR));

	always begin

	//0
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//1
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//2
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//3
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//4
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//5
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//6
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//7
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//8
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//9
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//10
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//11
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//12
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//13
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//14
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//15
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//16
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//17
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//18
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//19
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//20
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//21
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//22
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//23
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//24
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//25
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//26
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//27
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//28
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//29
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//30
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//31
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//32
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//33
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//34
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//35
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//36
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//37
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//38
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//39
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//40
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//41
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//42
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//43
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//44
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//45
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//46
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//47
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//48
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//49
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//50
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//51
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//52
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//53
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//54
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//55
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//56
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//57
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//58
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//59
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//60
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//61
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//62
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//63
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//64
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//65
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//66
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//67
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//68
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//69
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//70
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//71
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//72
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//73
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//74
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//75
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//76
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//77
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//78
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//79
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//80
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//81
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//82
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//83
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//84
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//85
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//86
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//87
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//88
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//89
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//90
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//91
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//92
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//93
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//94
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//95
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//96
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//97
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//98
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//99
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//100
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//101
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//102
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//103
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//104
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//105
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//106
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//107
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//108
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//109
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//110
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//111
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//112
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//113
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//114
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//115
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//116
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//117
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//118
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//119
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//120
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//121
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//122
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//123
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//124
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//125
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//126
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//127
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//128
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//129
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//130
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//131
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//132
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//133
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//134
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//135
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//136
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//137
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//138
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//139
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//140
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//141
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//142
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//143
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//144
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//145
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//146
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//147
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//148
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//149
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//150
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//151
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//152
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//153
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//154
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//155
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//156
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//157
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//158
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//159
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//160
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//161
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//162
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//163
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//164
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//165
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//166
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//167
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//168
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//169
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//170
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//171
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//172
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//173
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//174
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//175
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//176
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//177
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//178
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//179
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//180
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//181
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//182
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//183
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//184
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//185
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//186
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//187
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//188
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//189
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//190
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//191
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//192
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//193
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//194
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//195
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//196
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//197
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//198
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//199
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//200
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//201
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//202
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//203
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//204
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//205
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//206
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//207
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//208
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//209
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//210
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//211
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//212
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//213
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//214
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//215
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//216
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//217
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//218
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//219
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//220
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//221
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//222
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//223
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//224
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//225
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//226
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//227
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//228
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//229
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//230
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//231
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//232
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//233
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//234
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//235
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//236
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//237
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//238
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//239
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//240
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//241
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//242
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//243
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//244
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//245
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//246
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//247
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//248
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//249
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//250
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//251
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//252
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//253
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//254
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//255
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//256
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//257
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//258
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//259
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//260
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//261
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//262
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//263
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//264
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//265
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//266
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//267
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//268
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//269
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//270
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//271
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//272
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//273
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//274
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//275
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//276
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//277
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//278
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//279
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//280
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//281
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//282
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//283
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//284
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//285
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//286
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//287
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//288
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//289
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//290
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//291
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//292
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//293
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//294
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//295
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//296
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//297
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//298
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//299
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//300
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//301
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//302
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//303
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//304
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//305
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//306
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//307
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//308
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//309
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//310
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//311
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//312
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//313
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//314
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//315
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//316
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//317
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//318
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//319
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//320
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//321
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//322
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//323
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//324
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//325
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//326
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//327
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//328
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//329
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//330
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//331
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//332
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//333
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//334
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//335
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//336
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//337
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//338
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//339
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//340
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//341
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//342
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//343
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//344
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//345
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//346
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//347
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//348
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//349
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//350
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//351
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//352
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//353
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//354
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//355
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//356
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//357
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//358
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//359
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//360
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//361
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//362
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//363
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//364
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//365
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//366
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//367
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//368
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//369
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//370
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//371
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//372
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//373
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//374
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//375
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//376
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//377
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//378
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//379
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//380
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//381
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//382
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//383
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//384
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//385
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//386
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//387
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//388
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//389
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//390
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//391
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//392
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//393
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//394
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//395
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//396
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//397
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//398
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//399
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//400
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//401
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//402
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//403
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//404
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//405
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//406
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//407
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//408
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//409
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//410
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//411
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//412
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//413
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//414
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//415
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//416
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//417
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//418
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//419
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//420
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//421
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//422
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//423
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//424
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//425
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//426
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//427
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//428
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//429
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//430
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//431
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//432
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//433
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//434
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//435
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//436
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//437
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//438
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//439
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//440
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//441
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//442
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//443
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//444
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//445
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//446
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//447
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//448
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//449
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//450
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//451
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//452
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//453
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//454
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//455
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//456
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//457
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//458
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//459
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//460
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//461
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//462
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//463
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//464
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//465
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//466
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//467
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//468
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//469
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//470
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//471
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//472
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//473
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//474
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//475
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//476
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//477
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//478
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//479
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//480
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//481
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//482
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//483
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//484
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//485
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//486
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//487
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//488
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//489
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//490
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//491
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//492
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//493
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//494
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//495
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//496
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//497
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//498
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//499
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//500
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//501
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//502
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//503
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//504
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//505
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//506
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//507
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//508
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//509
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//510
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//511
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//512
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//513
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//514
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//515
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//516
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//517
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//518
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//519
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//520
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//521
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//522
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//523
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//524
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//525
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//526
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//527
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//528
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//529
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//530
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//531
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//532
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//533
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//534
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//535
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//536
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//537
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//538
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//539
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//540
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//541
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//542
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//543
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//544
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//545
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//546
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//547
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//548
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//549
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//550
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//551
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//552
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//553
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//554
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//555
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//556
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//557
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//558
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//559
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//560
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//561
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//562
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//563
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//564
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//565
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//566
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//567
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//568
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//569
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//570
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//571
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//572
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//573
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//574
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//575
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//576
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//577
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//578
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//579
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//580
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//581
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//582
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//583
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//584
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//585
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//586
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//587
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//588
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//589
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//590
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//591
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//592
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//593
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//594
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//595
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//596
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//597
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//598
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//599
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//600
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//601
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//602
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//603
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//604
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//605
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//606
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//607
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//608
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//609
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//610
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//611
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//612
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//613
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//614
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//615
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//616
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//617
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//618
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//619
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//620
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//621
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//622
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//623
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//624
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//625
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//626
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//627
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//628
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//629
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//630
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//631
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//632
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//633
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//634
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//635
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//636
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//637
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//638
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//639
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//640
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//641
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//642
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//643
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//644
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//645
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//646
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//647
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//648
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//649
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//650
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//651
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//652
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//653
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//654
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//655
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//656
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//657
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//658
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//659
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//660
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//661
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//662
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//663
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//664
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//665
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//666
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//667
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//668
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//669
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//670
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//671
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//672
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//673
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//674
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//675
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//676
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//677
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//678
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//679
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//680
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//681
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//682
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//683
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//684
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//685
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//686
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//687
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//688
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//689
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//690
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//691
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//692
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//693
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//694
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//695
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//696
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//697
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//698
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//699
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//700
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//701
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//702
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//703
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//704
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//705
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//706
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//707
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//708
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//709
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//710
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//711
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//712
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//713
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//714
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//715
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//716
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//717
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//718
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//719
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//720
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//721
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//722
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//723
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//724
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//725
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//726
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//727
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//728
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//729
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//730
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//731
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//732
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//733
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//734
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//735
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//736
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//737
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//738
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//739
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//740
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//741
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//742
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//743
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//744
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//745
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//746
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//747
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//748
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//749
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//750
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//751
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//752
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//753
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//754
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//755
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//756
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//757
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//758
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//759
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//760
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//761
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//762
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//763
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//764
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//765
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//766
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//767
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b0;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//768
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//769
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//770
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//771
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//772
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//773
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//774
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//775
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//776
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//777
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//778
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//779
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//780
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//781
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//782
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//783
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//784
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//785
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//786
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//787
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//788
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//789
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//790
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//791
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//792
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//793
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//794
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//795
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//796
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//797
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//798
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//799
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//800
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//801
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//802
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//803
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//804
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//805
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//806
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//807
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//808
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//809
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//810
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//811
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//812
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//813
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//814
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//815
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//816
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//817
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//818
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//819
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//820
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//821
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//822
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//823
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//824
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//825
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//826
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//827
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//828
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//829
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//830
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//831
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//832
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//833
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//834
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//835
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//836
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//837
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//838
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//839
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//840
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//841
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//842
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//843
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//844
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//845
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//846
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//847
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//848
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//849
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//850
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//851
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//852
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//853
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//854
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//855
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//856
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//857
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//858
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//859
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//860
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//861
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//862
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//863
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//864
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//865
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//866
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//867
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//868
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//869
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//870
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//871
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//872
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//873
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//874
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//875
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//876
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//877
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//878
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//879
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//880
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//881
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//882
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//883
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//884
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//885
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//886
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//887
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//888
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//889
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//890
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//891
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//892
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//893
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//894
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//895
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b0;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//896
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//897
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//898
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//899
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//900
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//901
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//902
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//903
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//904
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//905
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//906
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//907
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//908
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//909
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//910
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//911
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//912
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//913
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//914
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//915
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//916
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//917
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//918
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//919
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//920
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//921
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//922
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//923
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//924
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//925
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//926
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//927
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//928
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//929
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//930
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//931
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//932
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//933
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//934
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//935
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//936
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//937
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//938
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//939
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//940
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//941
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//942
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//943
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//944
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//945
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//946
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//947
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//948
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//949
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//950
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//951
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//952
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//953
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//954
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//955
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//956
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//957
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//958
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//959
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b0;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//960
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//961
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//962
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//963
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//964
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//965
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//966
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//967
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//968
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//969
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//970
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//971
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//972
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//973
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//974
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//975
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//976
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//977
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//978
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//979
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//980
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//981
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//982
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//983
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//984
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//985
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//986
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//987
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//988
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//989
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//990
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//991
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b0;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//992
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//993
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//994
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//995
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//996
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//997
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//998
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//999
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//1000
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//1001
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//1002
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//1003
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//1004
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//1005
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//1006
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//1007
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b0;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//1008
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//1009
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//1010
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//1011
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//1012
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//1013
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//1014
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//1015
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b0;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//1016
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//1017
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//1018
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//1019
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b0;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;

	//1020
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b0;

	//1021
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b0;
		TB_A[0] = 1'b1;

	//1022
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b0;

	//1023
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_EN = 1'b1;
	#5 clk = 1'b1;
	#5 TB_EN = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	#10 clk = 1'b0;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;


	#10 clk = 1'b1;
		TB_RST = 1'b1;
		TB_B[3] = 1'b1;
		TB_B[2] = 1'b1;
		TB_B[1] = 1'b1;
		TB_B[0] = 1'b1;
		TB_A[3] = 1'b1;
		TB_A[2] = 1'b1;
		TB_A[1] = 1'b1;
		TB_A[0] = 1'b1;
	end

endmodule